//----------------------------------------------------------------------
//                   Mentor Graphics Corporation
//----------------------------------------------------------------------
// Project         : divisor
// Unit            : vsequence4
// File            : vsequence4.svh
//----------------------------------------------------------------------
// Created by      : rgadea
// Creation Date   : 2022/05/23
//----------------------------------------------------------------------
// Title: 
//
// Summary:
//
// Description:
//
//----------------------------------------------------------------------

//----------------------------------------------------------------------
// vsequence4
//----------------------------------------------------------------------
class vsequence4 extends virtual_sequence_base;

  // factory registration macro
  `uvm_object_utils(vsequence4)

  //--------------------------------------------------------------------
  // new
  //--------------------------------------------------------------------   
  function new(string name = "vsequence4");
    super.new(name);
  endfunction: new

  //--------------------------------------------------------------------
  // body
  //--------------------------------------------------------------------   
  task body();
    sequence4 seq_a = sequence4::type_id::create("seq_a");
    seq_a.start(m_agente_unico_sequencer);
  endtask: body

endclass: vsequence4

