//----------------------------------------------------------------------
//                   Mentor Graphics Corporation
//----------------------------------------------------------------------
// Project         : divisor
// Unit            : vsequence3
// File            : vsequence3.svh
//----------------------------------------------------------------------
// Created by      : rgadea
// Creation Date   : 2022/05/23
//----------------------------------------------------------------------
// Title: 
//
// Summary:
//
// Description:
//
//----------------------------------------------------------------------

//----------------------------------------------------------------------
// vsequence3
//----------------------------------------------------------------------
class vsequence3 extends virtual_sequence_base;

  // factory registration macro
  `uvm_object_utils(vsequence3)

  //--------------------------------------------------------------------
  // new
  //--------------------------------------------------------------------   
  function new(string name = "vsequence3");
    super.new(name);
  endfunction: new

  //--------------------------------------------------------------------
  // body
  //--------------------------------------------------------------------   
  task body();
    sequence3 seq_a = sequence3::type_id::create("seq_a");
    seq_a.start(m_agente_unico_sequencer);
  endtask: body

endclass: vsequence3

